module slot(
input clk,
input rst,
input [1:0]status,
output [3:0] value

);
endmodule