module miniALU
(
	input wire in,
	output wire out
);

endmodule