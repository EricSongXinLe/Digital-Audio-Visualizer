module miniALU_top
(
	input [9:0] in,
	output [9:0] out
);
assign out = in;
endmodule